// @top: test_compact
// @category: test
// @compact: true

module test_compact(input [7:0] a, b, output [7:0] o);
    assign o = a & b;
endmodule
