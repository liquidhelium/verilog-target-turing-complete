// @top: basic_and
// @category: basic
module basic_and(input wire a, input wire b, output wire y);
  assign y = a & b;
endmodule
