// @top: basic_wire
// @category: basic
module basic_wire(input wire a, output wire y);
  assign y = a;
endmodule
