// @top: basic_or
// @category: basic
module basic_or(input wire a, input wire b, output wire y);
  assign y = a | b;
endmodule
