// @top: test_add
// @category: test
module test_add (
    input [7:0] a,
    input [7:0] b,
    output [7:0] y
);
    assign y = a + b;
endmodule
