// @top: bus_odd_31
// @category: new
module bus_odd_31(input wire [30:0] a, input wire [30:0] b, output wire [30:0] y);
  assign y = a & b;
endmodule
