// @top: const_test
// @category: const
module const_test(output wire [31:0] y);
    assign y = 32'hDEADBEEF;
endmodule
