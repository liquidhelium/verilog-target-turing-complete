// @top: basic_not
// @category: basic
module basic_not(input wire a, output wire y);
  assign y = ~a;
endmodule
